LIBRARY ieee;
use ieee.std_logic_1164.all;
use work.MIPS_components.all;

--16bit ALU
Entity ALU16 IS
	PORT (A,B: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			SEL: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			COUT,OVERFLOW,ZERO: OUT STD_LOGIC;
			F: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ALU16;

ARCHITECTURE Behavior of ALU16 IS
	SIGNAL SETsig,COUT1,COUT2,COUT3,ZERO0,ZERO1,ZERO2,ZERO3, DNC: STD_LOGIC;
	
BEGIN 
	ALULOW: 	  ALU4 PORT MAP(A(3 DOWNTO 0),  B(3 DOWNTO 0),  SETsig,SEL(2),SEL,COUT1,DNC,DNC,  ZERO0,F(3 DOWNTO 0));	--PORTMAP all of the ALUS
	ALULOWMED: ALU4 PORT MAP(A(7 DOWNTO 4),  B(7 DOWNTO 4),  '0',COUT1,SEL,COUT2,DNC,DNC,      ZERO1,F(7 DOWNTO 4));
	ALUHIGHMED:ALU4 PORT MAP(A(11 DOWNTO 8), B(11 DOWNTO 8), '0',COUT2,SEL,COUT3,DNC,DNC,      ZERO2,F(11 DOWNTO 8));
	ALUHIGH:   ALU4 PORT MAP(A(15 DOWNTO 12),B(15 DOWNTO 12),'0',COUT3,SEL,COUT,OVERFLOW,SETsig, ZERO3,F(15 DOWNTO 12));
	ZERO<= (ZERO0 AND ZERO1 AND ZERO2 AND ZERO3);

	
	

	
	

END Behavior;