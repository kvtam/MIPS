LIBRARY ieee;
use ieee.std_logic_1164.all;
use work.MIPS_components.all;



--16bit Adder
Entity ADD16 IS
	PORT(A,B :IN STD_LOGIC_VECTOR(15 DOWNTO 0);
         Cin :IN STD_LOGIC;
         S   :OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
         Cout:OUT  STD_LOGIC);
END ADD16;

ARCHITECTURE Behavior of ADD16 IS
	SIGNAL COUT0, COUT1, COUT2: STD_LOGIC;
	
BEGIN 
	ADD0: ADD4 PORT MAP(A(3 DOWNTO 0), B(3 DOWNTO 0), Cin,S(3 DOWNTO 0), COUT0);
	ADD1: ADD4 PORT MAP(A(7 DOWNTO 4), B(7 DOWNTO 4), COUT0,S(7 DOWNTO 4), COUT1);
	ADD2: ADD4 PORT MAP(A(11 DOWNTO 8), B(11 DOWNTO 8), COUT1,S(11 DOWNTO 8), COUT2);
	ADD3: ADD4 PORT MAP(A(15 DOWNTO 12), B(15 DOWNTO 12), COUT2,S(15 DOWNTO 12), COUT);
	
	
	
END Behavior;