LIBRARY ieee;
use ieee.std_logic_1164.all;
use work.MIPS_components.all;
--16bit 8 to 1 mux
Entity MUX8x16 IS
	PORT (D0,D1,D2,D3,D4,D5,D6,D7: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			s:	IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			Q: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END MUX8x16;

ARCHITECTURE Behavior of MUX8x16 IS

--	COMPONENT MUX4x4
--		PORT (D0,D1,D2,D3: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
--			s:	IN STD_LOGIC_VECTOR (1 DOWNTO 0);
--			Q: OUT STD_LOGIC_VECTOR (3 DOWNTO 0));
--	END COMPONENT;
	signal LOWBITS, HIGHBITS: STD_LOGIC_VECTOR(15 DOWNTO 0);
	BEGIN 
		
		
	low_bits_12to15: MUX4x4 PORT MAP (D0(15 DOWNTO 12), D1(15 DOWNTO 12), D2( 15 DOWNTO 12), D3(15 DOWNTO 12), s(1 DOWNTO 0), LOWBITS(15 DOWNTO 12));
	low_bits_8to11: MUX4x4 PORT MAP (D0(11 DOWNTO 8), D1(11 DOWNTO 8), D2( 11 DOWNTO 8), D3(11 DOWNTO 8), s(1 DOWNTO 0), LOWBITS(11 DOWNTO 8));
	low_bits_4to7: MUX4x4 PORT MAP (D0(7 DOWNTO 4), D1(7 DOWNTO 4), D2( 7 DOWNTO 4), D3(7 DOWNTO 4), s(1 DOWNTO 0), LOWBITS(7 DOWNTO 4));
	low_bits_0to3: MUX4x4 PORT MAP (D0(3 DOWNTO 0), D1(3 DOWNTO 0), D2( 3 DOWNTO 0), D3(3 DOWNTO 0), s(1 DOWNTO 0), LOWBITS(3 DOWNTO 0));
	
	high_bits_12to15: MUX4x4 PORT MAP (D4(15 DOWNTO 12), D5(15 DOWNTO 12), D6( 15 DOWNTO 12), D7(15 DOWNTO 12), s(1 DOWNTO 0), HIGHBITS(15 DOWNTO 12));
	high_bits_8to11: MUX4x4 PORT MAP (D4(11 DOWNTO 8), D5(11 DOWNTO 8), D6( 11 DOWNTO 8), D7(11 DOWNTO 8), s(1 DOWNTO 0), HIGHBITS(11 DOWNTO 8));
	high_bits_4to7: MUX4x4 PORT MAP (D4(7 DOWNTO 4), D5(7 DOWNTO 4), D6( 7 DOWNTO 4), D7(7 DOWNTO 4), s(1 DOWNTO 0), HIGHBITS(7 DOWNTO 4));
	high_bits_0to3: MUX4x4 PORT MAP (D4(3 DOWNTO 0), D5(3 DOWNTO 0), D6( 3 DOWNTO 0), D7(3 DOWNTO 0), s(1 DOWNTO 0), HIGHBITS(3 DOWNTO 0));
	
	with s(2) select
	Q<= LOWBITS when '0',
	HIGHBITS when '1';
	
END Behavior;
				