LIBRARY ieee;
use ieee.std_logic_1164.all;
use work.MIPS_components.all;

--4x16 dec
Entity DCD4x16 IS
	PORT (D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			EN:IN STD_LOGIC;
			Q: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END DCD4x16;

ARCHITECTURE Behavior of DCD4x16 IS
		Signal RES: STD_LOGIC_VECTOR(15 DOWNTO 0);
	BEGIN 
		LOWBITS: DCD3x8 PORT MAP(D(2 DOWNTO 0),(NOT D(3)),RES(7 DOWNTO 0));
		HIGHBITS: DCD3x8 PORT MAP(D(2 DOWNTO 0),D(3),RES(15 DOWNTO 8));
		WITH EN SELECT
			Q<="0000000000000000" WHEN '0',
			RES WHEN '1';
	
		
END Behavior;
				